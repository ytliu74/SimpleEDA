My Testbench

R1 node_1 node_2 1k
C1 node_2 node_3 1p
c1 node_3 node_1 1m

Ix gnd node_2 10

.print V(node_2)

.end