Test tran

V1 1 0 10
R1 1 2 1
L1 1 2 1
C1 2 0 1

.tran 1 10
.END