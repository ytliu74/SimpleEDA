A test for diode

R1 0 1 1
D1 2 0 d_model
V1 1 0 5

.end