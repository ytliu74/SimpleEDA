My Testbench

R1 node_1 node_2 1k
C1 node_2 node_3 1p
L1 node_3 node_1 1m

VIN node_2 node_1 4

.print V(node_2)

.end