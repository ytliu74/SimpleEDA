Test tran

V1 1 0 10
R1 1 2 1k
R2 2 0 4k

.dc V1 0 10 1
.END